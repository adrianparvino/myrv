module furbi(
    input clk_i,
    output [15:0] adr_o,
    input [31:0] dat_i,
    output [31:0] dat_o,
    output we_o,
    output sel_o,
    output stb_o,
    input ack_i,
    output cyc_o
);

furv furv()

endmodule
