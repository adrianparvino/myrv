module myrv(
  input program, 
  output reg pc
);

  

endmodule
